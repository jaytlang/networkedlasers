parameter EIDLE = 0;
parameter ENOV4 = 1;
parameter ESHDR = 2;
parameter EDEAD = 3;
parameter EPROT = 4;
parameter EFRAG = 5;
parameter EPDST = 6;
parameter EETYP = 7;
parameter ECSUM = 8;
parameter EPORT = 9;
parameter EGOOD = 'hffff;
parameter EARPQ = 'hff01;
parameter EECHO = 'hff02;
